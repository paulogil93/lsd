-- Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, the Altera Quartus Prime License Agreement,
-- the Altera MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Altera and sold by Altera or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- Generated by Quartus Prime Version 15.1.2 Build 193 02/01/2016 SJ Lite Edition
-- Created on Wed May 18 14:59:18 2016

LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY DrinksFSM IS
    PORT (
        clk : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        Vin : IN STD_LOGIC := '0';
        Cin : IN STD_LOGIC := '0';
        drink : OUT STD_LOGIC;
		  count : OUT STD_LOGIC_VECTOR(3 downto 0)
    );
END DrinksFSM;

ARCHITECTURE BEHAVIOR OF DrinksFSM IS
    TYPE type_fstate IS (S0,S1,S2,S3,S4,S5);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
	 SIGNAL s_count : unsigned(3 downto 0);
BEGIN
    PROCESS (clk,reg_fstate)
    BEGIN
        IF (clk='1' AND clk'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,Vin,Cin)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= S0;
            drink <= '0';
				s_count <= (others => '0');
        ELSE
            drink <= '0';
            CASE fstate IS
                WHEN S0 =>
						  s_count <= (others => '0');
                    IF (((Vin = '1') AND NOT((Cin = '1')))) THEN
                        reg_fstate <= S1;
								s_count <= s_count + 2;
                    ELSIF (((Cin = '1') AND NOT((Vin = '1')))) THEN
                        reg_fstate <= S3;
								s_count <= s_count + 5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S0;
                    END IF;

                    drink <= '0';
                WHEN S1 =>
                    IF (((Vin = '1') AND NOT((Cin = '1')))) THEN
                        reg_fstate <= S2;
								s_count <= s_count + 2;
                    ELSIF (((Cin = '1') AND NOT((Vin = '1')))) THEN
                        reg_fstate <= S4;
								s_count <= s_count + 5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S0;
                    END IF;

                    drink <= '0';
                WHEN S2 =>
                    IF (((Vin = '1') AND NOT((Cin = '1')))) THEN
                        reg_fstate <= S3;
								s_count <= s_count + 2;
                    ELSIF (((Cin = '1') AND NOT((Vin = '1')))) THEN
                        reg_fstate <= S5;
								s_count <= s_count + 5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S0;
                    END IF;

                    drink <= '0';
                WHEN S3 =>
                    IF (((Vin = '1') AND NOT((Cin = '1')))) THEN
                        reg_fstate <= S4;
								s_count <= s_count + 2;
                    ELSIF (((Cin = '1') AND NOT((Vin = '1')))) THEN
                        reg_fstate <= S5;
								s_count <= s_count + 5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S0;
                    END IF;

                    drink <= '0';
                WHEN S4 =>
                    IF (((Vin = '1') OR (Cin = '1'))) THEN
                        reg_fstate <= S5;
								IF(Vin = '1') THEN
									s_count <= s_count + 2;
								ELSIF(Cin = '1') THEN
									s_count <= s_count + 5;
								END IF;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S0;
                    END IF;

                    drink <= '0';
                WHEN S5 =>
                    reg_fstate <= S0;
                    drink <= '1';
                WHEN OTHERS => 
                    drink <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
	 
	 count <= std_logic_vector(s_count);
END BEHAVIOR;
